* C:\Users\91766\Desktop\sky130\serilizer\serilizer.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/08/22 20:53:50

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ Din Din_bar dac_bridge_2		
U7  Net-_U2-Pad8_ Net-_U10-Pad1_ Net-_U10-Pad2_ buffer		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ mux4to1		
U5  s1 s0 en0 Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ adc_bridge_3		
U4  data3 data2 data1 data0 Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ adc_bridge_4		
v1  data3 GND pulse		
v3  data1 GND pulse		
v5  s1 GND pulse		
v7  en0 GND pulse		
v6  s0 GND pulse		
U3  data3 plot_v1		
U1  data1 plot_v1		
U6  s1 plot_v1		
U8  s0 plot_v1		
U9  en0 plot_v1		
U11  Din plot_v1		
U12  Din_bar plot_v1		
X1  vdd Din Din_bar vbias voa vob vocm LVDR		
vdd1  vdd GND DC		
vbais1  vbias GND DC		
U15  voa plot_v1		
U17  vocm plot_v1		
U16  vob plot_v1		
v2  data2 GND pulse		
U13  data2 plot_v1		
v4  data0 GND pulse		
U14  data0 plot_v1		
scmode1  SKY130mode		

.end
